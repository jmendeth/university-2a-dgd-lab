library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;

entity CA2_BCD_8B is
  port ( Ca2 : in std_logic_vector(4 downto 0);
         BCD : out std_logic_vector(7 downto 0) );
end;

architecture logic of CA2_BCD_8B is
begin
end logic;